

<!DOCTYPE html>


<html lang="sv" class="no-js" dir="ltr">
<head about=" ">
    <meta charset="utf-8">
    <title></title>
    <meta name="viewport" content="width=device-width, initial-scale=1.0">
    <meta name="description" content="">
    <meta name="author" content="">
    <meta http-equiv="Content-Type" content="application/xhtml+xml; charset=utf-8" />
    <meta name="keywords" content="">
    <link rel="stylesheet" href="https://cdn.jsdelivr.net/npm/bulma@0.9.0/css/bulma.min.css">
    <link rel="stylesheet" href="https://cdn.jsdelivr.net/npm/@creativecommons/vocabulary/css/vocabulary.css">
</head>
<body typeoff="cc:License">
  <style>svg { height: 73px; }</style>

<header>
  <nav class="navbar">
    <div class="navbar-brand">
      <a id="cc-logo" class="has-text-black" href="https://creativecommons.org" rel="home">
        <svg
          xmlns="http://www.w3.org/2000/svg"
          preserveAspectRatio="xMidYMid meet"
          viewBox="0 0 304 73">
        <!-- Automatically finds ID amongst all assets loaded using `patchAssetIntoDom()` -->
          <use href="#logomark"></use>
        </svg>
      </a>
      <a role="button" class="navbar-burger is-active" aria-label="menu" aria-expanded="false">
        <span aria-hidden="true"></span>
        <span aria-hidden="true"></span>
        <span aria-hidden="true"></span>
      </a>
    </div>
    <div class="navbar-menu is-active">
      <div class="navbar-end">
        <div class="navbar-item has-dropdown is-hoverable">
          <a class="navbar-link is-arrowless">Who We Are<i class="icon caret-down"></i></a>
          <div class="navbar-dropdown">
            <a class="navbar-item">Item 1</a>
            <a class="navbar-item">Item 2</a>
            <a class="navbar-item">Item 3</a>
          </div>
        </div>
        <div class="navbar-item has-dropdown is-hoverable">
          <a class="navbar-link is-arrowless">What We Do<i class="icon caret-down"></i></a>
          <div class="navbar-dropdown">
            <a class="navbar-item">Item 1</a>
            <a class="navbar-item">Item 2</a>
            <a class="navbar-item">Item 3</a>
          </div>
        </div>
        <a class="navbar-item">
          Our Impact<i class="icon external-link"></i>
        </a>
        <a class="navbar-item">
          News
        </a>
      </div>
    </div>
  </nav>
</header>

<style>
  html[dir="rtl"] .has-dropdown .navbar-link {
      flex-direction: row-reverse;
  }

  html[dir="rtl"] .navbar-end {
      margin-right: auto;
      margin-left: 0;
      justify-content: flex-start;
  }
</style>

  <main>
    <div class="level padding-left-big padding-right-large padding-vertical-normal">
          


<a class="skip-link" href="#content" >Hoppa över till innehåll</a>

<style>
  a.skip-link {
    left:-999px;
    position:absolute;
    top:auto;
    width:1px;
    height:1px;
    overflow:hidden;
    z-index:-999;
}
a.skip-link:focus, a.skip-link:active {
    color: black;
    font-weight: bolder;
    left: auto;
    top: auto;
    width: 30%;
    height: auto;
    overflow:auto;
    margin: 10px 35%;
    padding:5px;
    background-color: rgb(255, 255, 255);
    border-top: 10px solid rgb(60, 92, 153);
    border-bottom: 5px solid rgb(176, 176, 176);
    border-left: 5px solid rgb(176, 176, 176);
    border-right: 5px solid rgb(176, 176, 176);
    text-align:center;
    font-size:1.2em;
    z-index:999;
}
</style>

          <nav class="breadcrumb level-left caption bold" aria-label="breadcrumbs">
            <ul>
                <li><a href="/">Hem</a></li>
                <li><a href="/licenses/">Licenses</a></li>
                
  <li class="is-active"><a href="/licenses/by-sa/4.0/legalcode.sv" aria-current="page displayed">Legal Code for CC BY-SA 4.0</a></li>

            </ul>
          </nav>
          
            


<div class="locale level-right level-item has-text-black" >
  Languages available
  <div class="control margin-left-small">
    <div class="select">
      <select id="languages-dropdown">
        
        <option disabled>Select</option>

        
          <option
            id="option-id"
            
            value="id"
            data-link="/licenses/by-sa/4.0/legalcode.id"
          >
            Bahasa Indonesia
          </option>
        
          <option
            id="option-eu"
            
            value="eu"
            data-link="/licenses/by-sa/4.0/legalcode.eu"
          >
            Basque
          </option>
        
          <option
            id="option-de"
            
            value="de"
            data-link="/licenses/by-sa/4.0/legalcode.de"
          >
            Deutsch
          </option>
        
          <option
            id="option-en"
            
            value="en"
            data-link="/licenses/by-sa/4.0/legalcode"
          >
            English
          </option>
        
          <option
            id="option-es"
            
            value="es"
            data-link="/licenses/by-sa/4.0/legalcode.es"
          >
            español
          </option>
        
          <option
            id="option-fr"
            
            value="fr"
            data-link="/licenses/by-sa/4.0/legalcode.fr"
          >
            français
          </option>
        
          <option
            id="option-hr"
            
            value="hr"
            data-link="/licenses/by-sa/4.0/legalcode.hr"
          >
            Hrvatski
          </option>
        
          <option
            id="option-it"
            
            value="it"
            data-link="/licenses/by-sa/4.0/legalcode.it"
          >
            italiano
          </option>
        
          <option
            id="option-lv"
            
            value="lv"
            data-link="/licenses/by-sa/4.0/legalcode.lv"
          >
            latviešu
          </option>
        
          <option
            id="option-lt"
            
            value="lt"
            data-link="/licenses/by-sa/4.0/legalcode.lt"
          >
            Lietuviškai
          </option>
        
          <option
            id="option-mi"
            
            value="mi"
            data-link="/licenses/by-sa/4.0/legalcode.mi"
          >
            Māori
          </option>
        
          <option
            id="option-nl"
            
            value="nl"
            data-link="/licenses/by-sa/4.0/legalcode.nl"
          >
            Nederlands
          </option>
        
          <option
            id="option-no"
            
            value="no"
            data-link="/licenses/by-sa/4.0/legalcode.no"
          >
            norsk
          </option>
        
          <option
            id="option-pl"
            
            value="pl"
            data-link="/licenses/by-sa/4.0/legalcode.pl"
          >
            polski
          </option>
        
          <option
            id="option-pt"
            
            value="pt"
            data-link="/licenses/by-sa/4.0/legalcode.pt"
          >
            Português
          </option>
        
          <option
            id="option-ro"
            
            value="ro"
            data-link="/licenses/by-sa/4.0/legalcode.ro"
          >
            Română
          </option>
        
          <option
            id="option-sl"
            
            value="sl"
            data-link="/licenses/by-sa/4.0/legalcode.sl"
          >
            Slovenščina
          </option>
        
          <option
            id="option-fi"
            
            value="fi"
            data-link="/licenses/by-sa/4.0/legalcode.fi"
          >
            suomi
          </option>
        
          <option
            id="option-sv"
            selected
            value="sv"
            data-link="/licenses/by-sa/4.0/legalcode.sv"
          >
            svenska
          </option>
        
          <option
            id="option-tr"
            
            value="tr"
            data-link="/licenses/by-sa/4.0/legalcode.tr"
          >
            Türkçe
          </option>
        
          <option
            id="option-cs"
            
            value="cs"
            data-link="/licenses/by-sa/4.0/legalcode.cs"
          >
            česky
          </option>
        
          <option
            id="option-el"
            
            value="el"
            data-link="/licenses/by-sa/4.0/legalcode.el"
          >
            Ελληνικά
          </option>
        
          <option
            id="option-ru"
            
            value="ru"
            data-link="/licenses/by-sa/4.0/legalcode.ru"
          >
            Русский
          </option>
        
          <option
            id="option-uk"
            
            value="uk"
            data-link="/licenses/by-sa/4.0/legalcode.uk"
          >
            Українська
          </option>
        
          <option
            id="option-ar"
            
            value="ar"
            data-link="/licenses/by-sa/4.0/legalcode.ar"
          >
            العربيّة
          </option>
        
          <option
            id="option-ja"
            
            value="ja"
            data-link="/licenses/by-sa/4.0/legalcode.ja"
          >
            日本語
          </option>
        
          <option
            id="option-zh-Hans"
            
            value="zh-Hans"
            data-link="/licenses/by-sa/4.0/legalcode.zh-Hans"
          >
            简体中文
          </option>
        
          <option
            id="option-zh-Hant"
            
            value="zh-Hant"
            data-link="/licenses/by-sa/4.0/legalcode.zh-Hant"
          >
            繁體中文
          </option>
        
          <option
            id="option-ko"
            
            value="ko"
            data-link="/licenses/by-sa/4.0/legalcode.ko"
          >
            한국어
          </option>
        

        
      </select>
    </div>
    <div class="icon is-small is-left">
      <!-- TODO Add icons here -->
    </div>
  </div>
</div>

<script>
  const select = document.getElementById("languages-dropdown")

  select.addEventListener("input", function () {
    const language_code = select.value
    const option = document.getElementById("option-" + language_code)
    window.location.href = option.dataset.link
  })
</script>

          
    </div>
    <section id="content" class="padding-horizontal-larger">
      
<div class="columns">
  <div class="column is-one-quarter"></div>
  <div class="column columns padding-vertical-normal">
    <div class="column is-three-quarters padding-top-normal">
      Version 4.0 &#8226;
      See the <a href="#">errata page</a> for any corrections and the date of change
      
    </div>
    <div class="column">
      <button id="next-btn" class="button tiny is-pulled-right" data-href="/licenses/by-sa/4.0/deed.sv">See the deed</button>
    </div>
  </div>
</div>

      
  <div class="columns">
    

<div class="column is-one-quarter sidebar-container">
  <aside class="menu sidebar-menu">
    <a class="link has-text-black is-block padding-bottom-normal" href="#legal-code-body">


Erkännande-DelaPåSammaVillkor 4.0 Internationell

</a>
    <ul class="menu-list" >
      <li>
        <ul>
          
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class="is-block column" href="#s1">Avsnitt 1 – Definitioner.</a>
          </li>
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class="is-block column" href="#s2">Avsnitt 2 – Omfattning.</a>
          </li>
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class="is-block column" href="#s3">Avsnitt 3 - Licensvillkor.</a>
          </li>
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class="is-block column" href="#s4">Avsnitt 4 – Sui Generis-rättigheter för Databaser.</a>
          </li>
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class="is-block column" href="#s5">Avsnitt 5 - Friskrivning från utfästelser och begränsning av ansvar.</a>
          </li>
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class=" is-block column" href="#s6">Avsnitt 6 – Giltighetstid och uppsägning.</a>
          </li>
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class="is-block column" href="#s7">Avsnitt 7 – Övriga villkor.</a>
          </li>
          <li class="columns">
            <div class="body-bigger is-inline-block column is-1 py-0 my-0">&#8226;</div>
            <a class=" is-block column" href="#s8">Avsnitt 8 – Tolkning.</a>
          </li>
        </ul>
      </li>
    </ul>
  </aside>
</div>

    <div class="column">
      



<div id="licenses-header" class="padding-larger margin-bottom-bigger has-text-black is-hidden-touch is-hidden-desktop-only" >
  <h2 class="is-vcentered">
    
      <span class="padding-right-bigger">
      
        





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


        





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


        





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


        





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      
      </span>

    CC BY-SA 4.0 
  </h2>
  
  <h1 class="b-header">


Erkännande-DelaPåSammaVillkor 4.0 Internationell

</h1>
</div>

<div id="licenses-header" class="padding-larger margin-bottom-bigger has-text-black is-hidden-widescreen" >
  <h2 class="has-text-centered">
    
      <span>
      
        





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


        





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


        





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


        





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-big padding-bottom-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      
      </span>
  </h2>
  <h2 class="has-text-centered is-hidden-touch is-hidden-desktop-only padding-left-normal">CC BY-SA 4.0</h2>
  <h3 class="has-text-centered is-hidden-touch">CC BY-SA 4.0</h3>
  <h4 class="has-text-centered is-hidden-desktop-only is-hidden-widescreen">CC BY-SA 4.0</h4>
  <h2 class="b-header has-text-centered">


Erkännande-DelaPåSammaVillkor 4.0 Internationell

</h2>
</div>

<style>
  #licenses-header {
    background-color: rgb(255, 255, 255);
    border-top: 10px solid rgb(60, 92, 153);
    border-bottom: 5px solid rgb(176, 176, 176);
    border-left: 5px solid rgb(176, 176, 176);
    border-right: 5px solid rgb(176, 176, 176);
  }
</style>

      



<div id="about-cc-and-license" class="padding-bigger has-background-info-light" >
  <h4 class="padding-bottom-normal is-vcentered b-header"><i class="info icon padding-right-normal"></i>About the license and Creative Commons</h4>
  <p class="has-text-black padding-left-big">
    Creative Commons Corporation ("Creative Commons") is not a law firm and does not provide legal services or legal advice. Distribution of Creative Commons public licenses does not create a lawyer-client or other relationship. Creative Commons makes its licenses and related information available on an "as-is" basis. Creative Commons gives no warranties regarding its licenses, any material licensed under their terms and conditions, or any related information. Creative Commons disclaims all liability for damages resulting from their use to the fullest extent possible.
  </p>
</div>

      


<div id="about-cc-and-license" class="padding-bigger margin-top-bigger has-background-info-light" >
  <h4 class="level is-vcentered b-header">Using Creative Commons Public Licenses</h4>
  <p class="has-text-black body-big">
    Creative Commons public licenses provide a standard set of terms and conditions that creators and other rights holders may use to share original works of authorship and other material subject to copyright and certain other rights specified in the public license below. The following considerations are for informational purposes only, are not exhaustive, and do not form part of our licenses.
  </p>
  <hr class="divider">
  <div>
    <h4 class="level is-vcentered b-header">Considerations for licensors<span class="level-right"><i class="angle-down icon" data-consideration="1" data-direction="down"><span class="is-sr-only">Show Considerations for Licensors</span></i></span></h4>
    <p class="has-text-black body-big is-hidden">
    Our public licenses are intended for use by those authorized to give the public permission to use material in ways otherwise restricted by copyright and certain other rights. Our licenses are irrevocable. Licensors should read and understand the terms and conditions of the license they choose before applying it. Licensors should also secure all rights necessary before applying our licenses so that the public can reuse the material as expected. Licensors should clearly mark any material not subject to the license. This includes other CC-licensed material, or material used under an exception or limitation to copyright. <a href="https://wiki.creativecommons.org/wiki/Considerations_for_licensors_and_licensees#Considerations_for_licensors">More considerations for licensors.</a>
    </p>
  </div>
  <hr class="divider">
  <div>
    <h4 class="level is-vcentered b-header">Considerations for the public<span class="level-right"><i class="angle-down icon" data-consideration="2" data-direction="down"><span class="is-sr-only">Show Considerations for the Public</span></i></span></h4>
    <p class="has-text-black body-big is-hidden">
    By using one of our public licenses, a licensor grants the public permission to use the licensed material under specified terms and conditions. If the licensor’s permission is not necessary for any reason–for example, because of any applicable exception or limitation to copyright–then that use is not regulated by the license. Our licenses grant only permissions under copyright and certain other rights that a licensor has authority to grant. Use of the licensed material may still be restricted for other reasons, including because others have copyright or other rights in the material. A licensor may make special requests, such as asking that all changes be marked or described. Although not required by our licenses, you are encouraged to respect those requests where reasonable. <a href="https://wiki.creativecommons.org/wiki/Considerations_for_licensors_and_licensees#Considerations_for_licensees">More considerations for the public.</a>
    </p>
  </div>
</div>

<style>
  [dir="rtl"] .has-background-info-light .divider {
      margin-right: -2rem;
  }
  [dir="ltr"] .has-background-info-light .divider {
      margin-left: -2rem;
  }

  .has-background-info-light .divider {
      width: calc(100% + 4rem);
      background-color: #b0b0b0;
  }
</style>

      
<div id="legal-code-body" class="padding-larger margin-top-bigger has-text-black">
  

<h3 class="is-vcentered is-hidden-touch">
  
    <span class="padding-right-bigger">
    
      





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


    </span>
  CC BY-SA 4.0
</h3>
<h3 class="is-vcentered is-hidden-desktop is-hidden-mobile has-text-centered">
  
    <span class="padding-right-big">
    
      





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


    </span>
    CC BY-SA 4.0
</h3>
<h3 class="is-hidden-tablet has-text-centered">
  
    <span>
    
      





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


      





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


      





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


      





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


    </span>
</h3>
<h4 class="has-text-centered is-hidden-tablet padding-left-normal">CC BY-SA 4.0</h4>
<h2 class="margin-bottom-larger b-header is-hidden-touch">


Erkännande-DelaPåSammaVillkor 4.0 Internationell

</h2>
<h3 class="margin-bottom-larger b-header is-hidden-desktop has-text-centered">


Erkännande-DelaPåSammaVillkor 4.0 Internationell

</h3>

  <div id="plain-text-marker"> 
    <h3 class="padding-bottom-normal b-header">
      
        Creative Commons Erkännande-DelaPåSammaVillkor 4.0 Internationell Publik Licens
      
    </h3>
    <p class="body-big padding-bottom-larger">
    
    Genom att nyttja Licensrättigheterna (definierade nedan), accepterar och godkänner Du att Du är bunden av villkoren i denna Creative Commons Erkännande-DelaPåSammaVillkor 4.0 Internationella Publika Licens ("Publik Licens"). I den mån den Publika Licensen kan tolkas som ett kontrakt, beviljas Du Licensrättigheterna under förutsättning att Du accepterar dessa villkor, och Licensgivaren beviljar Dig sådana rättigheter i förhållande till den nytta Licensgivaren har genom att göra Licensmaterialet tillgängligt under dessa villkor.
    
    </p>
    

    <!-- Section 1. Definitions. -->
    <div class="padding-bottom-larger">
      <p id="s1" class="body-bigger padding-bottom-normal"><strong>Avsnitt 1 – Definitioner.</strong></p>
      
      <ol type="a" class="body-big padding-left-normal">

          

          <li id="s1a_adapted_material" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Bearbetning</span> avses material som är föremål för Upphovsrätt eller Liknande Rättigheter som härrör från eller är baserat på Licensmaterialet och där Licensmaterialet har översatts, ändrats, arrangerats, omvandlats, eller på annat sätt modifierats på ett sätt som kräver tillstånd för Upphovsrätt eller Liknande Rättigheter som innehas av Licensgivaren. För tillämpningen av den här Publika Licensen har en Bearbetning alltid skapats när Licensmaterialet är synkroniserat med rörlig bild och utgör ett musikaliskt verk, ett framförande eller en ljudupptagning.</div>
          </li>

          
            <li id="s1b_adapters_license" class="padding-bottom-normal">
              <div class="padding-left-normal"><span style="text-decoration: underline;">Med Bearbetningslicens</span> avses den licens Du tillämpar rörande Din Upphovsrätt och och Liknande Rättigheter när du bidrar till en Bearbetning enligt villkoren i denna Publika Licens.</div>
            </li>
          

          

          
            <li id="s1c_by_sa_compatible_license" class="padding-bottom-normal">
              <div class="padding-left-normal"><span style="text-decoration: underline;"> Med BY-SA-Kompatibel Licens</span> avses en licens som har registrerats på <a href="//creativecommons.org/compatiblelicenses"> creativecommons.org/compatiblelicenses</a>, godkänd av Creative Commons som huvudsakligen jämförlig med denna Publika Licens.</div>
            </li>
          

          <li id="s1d_copyright_and_similar_rights" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Upphovsrätt eller Liknande Rättigheter</span> avses upphovsrätt och/eller liknande rättigheter närbesläktade med upphovsrätt, vilket utan begränsning inkluderar framförande, utsändning, ljudinspelning och Sui Generis-rättigheter för Databaser, oavsett hur rättigheterna är märkta eller kategoriserade. För tillämpningen av denna Publika Licens är de rättigheter som anges i avsnitt <a href="#s2b">2(b)(1)-(2)</a> inte Upphovsrätt eller Liknande Rättigheter.</div>
          </li>

          <li id="s1e_effective_technological_measures" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Tekniska Skyddsåtgärder</span> avses de åtgärder som inte utan behörighet får kringgås enligt de lagar som uppfyller skyldigheterna enligt artikel 11 i WIPO Copyright Treaty (WIPOs Upphovsrättsfördrag) som antogs den 20 december 1996 och/eller genom liknande internationella överenskommelser.</div>
          </li>

          <li id="s1f_exceptions_and_limitations" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Undantag och Begränsningar</span> avses "fair use", "fair dealing" och/eller varje annan form av undantag från eller inskränkningar i Upphovsrätt eller Liknande rättigheter som gäller för Din användning av Licensmaterialet.</div>
          </li>

          

          
            <li id="s1g_license_elements_sa" class="padding-bottom-normal">
              <div class="padding-left-normal"><span style="text-decoration: underline;">Med Grundlicens</span> avses de licensegenskaper som anges i rubriken till en Creative Commons Publik Licens. Grundlicenser för denna Publika Licens är ”Erkännande” och ”DelaPåSammaVillkor”.</div>
            </li>
          

          <li id="s1h_licensed_material" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Licensmaterialet</span> avses det konstnärliga eller litterära verk, databas, eller annat material som Licensgivaren tillämpat denna Publika Licens för.</div>
          </li>

          <li id="s1i_licensed_rights" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Licensrättigheter</span> avses de rättigheter som Du beviljas enligt villkoren i denna Publika Licens, vilka är begränsade till all Upphovsrätt eller Liknande rättigheter som gäller för Din användning av Licensmaterialet och som Licensgivaren har behörighet att licensiera.</div>
          </li>

          <li id="s1j_licensor" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Licensgivaren</span> avses den fysiska eller juridiska person som beviljar rättigheter enligt denna Publika Licens.</div>
          </li>

          

          <li id="s1k_share" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Dela</span> avses att tillhandahålla material till allmänheten på alla sätt och vis som kräver tillstånd enligt Licensrättigheterna, såsom mångfaldigande, offentlig visning, offentligt framförande, distribution, spridning, kommunikation, eller import, och att göra materialet tillgängligt för allmänheten även på de sätt som medlemmar av allmänheten kan få tillgång till material från en plats och vid en tidpunkt som de väljer själva.</div>
          </li>

          <li id="s1l_sui_generis_database_rights" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Sui Generis-rättigheter för Databaser</span> menas rättigheter vid sidan av upphovsrätt som följer av Europaparlamentets och rådets direktiv 96/9/EU av den 11 mars 1996 om rättsligt skydd för databaser, så som det är implementerat och/eller förändrat eller ersatt, liksom andra huvudsakligen likvärdiga rättigheter runtom i världen.</div>
          </li>

          <li id="s1m_you" class="padding-bottom-normal">
            <div class="padding-left-normal"><span style="text-decoration: underline;">Med Du</span> avses den fysiska eller juridiska person som utövar Licensrättigheterna enligt denna Publika Licens. Din, Ditt eller Dina har motsvarande betydelse. <strong>Dig</strong> har en liknande betydelse.</div>
          </li>
      </ol>
    </div>

    <!-- Section 2. Scope. -->
    <div class="padding-bottom-larger">
      <p id="s2" class="body-bigger padding-bottom-normal"><strong>Avsnitt 2 – Omfattning.</strong></p>
      <ol type="a" class="body-big padding-left-normal">
        <li id="s2a" class="padding-left-normal"><strong>Tillstånd enligt licens</strong>.
        <ol class="padding-left-normal padding-vertical-normal">
          <li id="s2a1" class="padding-left-normal padding-bottom-normal">Med förbehåll för villkoren i denna Publika Licens, beviljar Licenstagaren en global, royalty-fri, icke-vidarelicensierbar, icke-exklusiv och oåterkallelig rätt att nyttja Licensrättigheterna i Licensmaterialet till att:
            <ol type="A" class="padding-left-normal padding-vertical-normal">
            
              <li id="s2a1A" class="padding-left-normal padding-bottom-normal">mångfaldiga och Dela Licensmaterialet, helt eller delvis; och</li>
            

            
              <li id="s2a1B" class="padding-left-normal padding-bottom-small">skapa, mångfaldiga och Dela Bearbetningar.</li>
            

            </ol>
          </li>
          <li id="s2a2" class="padding-left-normal padding-bottom-normal"><strong>Undantag och Begränsningar</strong>. För att undvika osäkerhet: när Ditt nyttjande av ett verk omfattas av inskränkningar i lagen gäller inte denna Publika Licens, och Du behöver inte tillämpa licensensvillkoren.</li>
          <li id="s2a3" class="padding-left-normal padding-bottom-normal"><strong>Giltighetstiden</strong>. Giltighetstiden för denna Publika Licens anges i avsnitt <a href="#s6a">6(a)</a>.</li>
          <li id="s2a4" class="padding-left-normal padding-bottom-normal"><strong>Medieformer och format; tekniska ändringar tillåts</strong>. Licensgivaren ger Dig rätt att nyttja Licensrättigheterna i alla nu kända och kommande medieformer och format, och att vidta de tekniska anpassningar som krävs för det. Licensgivaren avstår från och/eller samtycker till att inte hävda någon rätt eller behörighet för att förbjuda Dig från att göra de nödvändiga tekniska anpassningar som krävs för att nyttja Licensieringsrättigheterna, däribland de tekniska anpassningar som krävs för att kringgå Tekniska skyddsåtgärder. Såvitt gäller tillämpningen av denna Publika Licens har Bearbetningar aldrig skapats genom anpassningar som är godkända enligt detta avsnitt <a href="#s2a4">2(a)(4)</a>.</li>
          <li id="s2a5" class="padding-left-normal padding-bottom-small">
            <span style="text-decoration: underline;">Senare nyttjare</span>.
            <div class="para">
              <ol type="A" class="padding-left-normal padding-vertical-normal">

                  

                  <li id="s2a5A_offer" class="padding-left-normal padding-bottom-normal"><span style="text-decoration: underline;">Erbjudande från Licensgivaren - Licensmaterialet</span>. Varje mottagare av Licensmaterialet får automatiskt ett erbjudande från Licensgivaren att nyttja de Licensrättigheterna enligt villkoren i denna Publika Licens.</li>

                  
                    <li id="s2a5B_adapted_material" class="padding-left-normal padding-bottom-normal"><span style="text-decoration: underline;">Tilläggserbjudande från Licensgivaren -- Bearbetningar</span>. Varje mottagare av Bearbetningar från Dig får automatiskt ett erbjudande från Licensgivaren att nyttja Licensrättigheterna som hör till Bearbetningen enligt villkoren i Bearbetningslicensen som Du tillämpar.</li>
                  

                  <li id="s2a5C_no_restrictions" class="padding-left-normal padding-bottom-small"><span style="text-decoration: underline;">Inga restriktioner för senare nyttjande</span>. Du får inte erbjuda eller införa något ytterligare eller annat villkor eller tillämpa någon Teknisk Skyddsåtgärd för Licensmaterialet om det innebär en begränsning av nyttjandet av Licensrättigheterna för någon mottagare av Licensmaterialet.</li>

              </ol>
            </div>
          </li>
          <li id="s2a6" class="padding-left-normal padding-bottom-small"><span style="text-decoration: underline;">Inget godkännande</span>. . Ingenting i denna Publika Licens utgör eller kan tolkas som tillstånd för att hävda eller antyda att Du eller Din användning av Licensmaterialet hör samman med eller är sponsrad, godkänd, eller beviljad officiell status av Licensgivaren eller andra som har rätt till erkännande enligt avsnitt <a href="#s3a1Ai">3(a)(1)(A)(i)</a>.</li>
        </ol>

        <li id="s2b" class="padding-left-normal"><strong>Andra rättigheter</strong>.
          <ol class="padding-left-normal padding-vertical-normal">
            <li id="s2b1" class="padding-left-normal padding-bottom-normal">Ideella rättigheter, såsom rätten till integritet, är inte licensierade under denna Publika Licens. Det gäller även publicitet, integritet, och/eller andra motsvarande personliga rättigheter; I den mån det är möjligt avstår dock Licensgivaren från och/eller samtycker till att inte hävda dylika rättigheter som hen innehar i den begränsade omfattning som krävs för att tillåta Dig att nyttja Licensrättigheterna, men inte i övrigt.</li>
            <li id="s2b2" class="padding-left-normal padding-bottom-normal">Patent och varumärkesrättigheter licensieras inte under denna Publika Licens.</li>
          
            <li id="s2b3" class="padding-left-normal padding-bottom-small">Licensgivaren avstår i möjligaste mån från rätten att erhålla royalty från Dig för nyttjandet av Licensrättigheterna, oavsett det sker direkt eller genom en upphovsrättsorganisation med stöd av ett frivilligt eller dispositivt lagstadgat eller obligatoriskt licenssystem. I alla andra fall förbehåller sig Licensgivaren uttryckligen rätten att erhålla sådan royalty.</li>
          
          </ol>
        </li>
      </ol>
    </div>

    <!-- Section 3. License Conditions. -->
    <div class="padding-bottom-larger">
      <p id="s3" class="body-bigger padding-bottom-normal"><strong>Avsnitt 3 - Licensvillkor.</strong></p>

      <p class="body-big padding-bottom-normal">Ditt nyttjande av Licensrättigheterna omfattas uttryckligen av följande villkor.</p>

      <ol type="a" class="body-big padding-left-normal">
        <li id="s3a" class="padding-left-normal padding-bottom-normal"><p><strong>Erkännande</strong>.</p>
          <ol type="1" class="padding-left-normal padding-vertical-normal">
            <li id="s3a1" class="padding-left-normal padding-bottom-normal">
              <p>Om Du Delar Licensmaterialet (inclusive i ändrad form), måste Du:</p>
              <ol type="A" class="padding-left-normal padding-vertical-normal">
                  <li id="s3a1A" class="padding-left-normal padding-bottom-small">behålla följande om det tillhandahålls av Licensgivaren tillsammans med Licensmaterialet:
                    <ol type="i" class="padding-left-normal padding-vertical-normal">
                        <li id="s3a1Ai" class="padding-left-normal padding-bottom-normal">identifiering av skaparen (-arna) av Licensmaterialet och andra som ska erkännas, på varje rimligt sätt som begärts av Licensgivaren (inbegripet pseudonym om sådan angivits);</li>
                        <li id="s3a1Aii" class="padding-left-normal padding-bottom-normal">ett meddelande om upphovsrätt;</li>
                        <li id="s3a1Aiii" class="padding-left-normal padding-bottom-normal">ett meddelande som hänvisar till denna Publika Licens;</li>
                        <li id="s3a1Aiv" class="padding-left-normal padding-bottom-normal">ett meddelande som hänvisar till friskrivning från garantier;</li>
                        <li id="s3a1Av" class="padding-left-normal padding-bottom-small">en URI eller hyperlänk till Licensmaterialet i den mån detta är rimligt genomförbart.</li>
                    </ol>
                  </li>
                  <li id="s3a1B" class="padding-left-normal padding-bottom-normal">ange om Du har ändrat i Licensmaterialet och bevara uppgifter om alla eventuella tidigare ändringar; och</li>
                  <li id="s3a1C" class="padding-left-normal padding-bottom-small">ange att Licensmaterialet är licensierat under denna Publika Licens och inkludera texten om, eller URI:en eller hyperlänken till, denna Publika Licens.</li>
              </ol>
            </li>
            <li id="s3a2" class="padding-left-normal padding-bottom-normal">Du kan uppfylla villkoren i avsnitt <a href="#s3a1">3(a)(1)</a> på varje rimligt sätt med tanke på det medium, sätt och sammanhang i vilket Du Delar Licensmaterialet. Till exempel kan det vara rimligt att uppfylla villkoren genom att tillhandahålla en URI eller hyperlänk till en resurs som innehåller den information som krävs.</li>
            
              <li id="s3a3" class="padding-left-normal padding-bottom-small">På begäran av Licensgivaren måste Du, i den mån det är rimligt genomförbart, avlägsna sådan information som krävs enligt avsnitt <a href="#s3a1A">3(a)(1)(A)</a>.</li>
              
            
          </ol>
        </li>

        
          <li id="s3b" class="padding-left-normal padding-bottom-normal"><strong>DelaPåSammaVillkor</strong>.
            <p class="padding-top-normal padding-bottom-normal">Om Du Delar de Bearbetningar Du har skapat gäller även följande villkor som tillägg till villkoren i avsnitt <a href="#s3a">3(a)</a>.</p>
            <ol class="padding-left-normal">
              <li id="s3b1" class="padding-left-normal padding-bottom-normal">Den Bearbetningslicens som Du tillämpar måste vara en Creative Commons-licens med samma typ av Grundlicens, i denna version eller senare, eller en BY-SA-kompatibel Licens.</li>
              <li id="s3b2" class="padding-left-normal padding-bottom-normal">Du måste inkludera texten om, eller URI:en eller hyperlänken till den Bearbetningslicens som Du tillämpar. Du kan uppfylla detta villkor på varje rimligt sätt med tanke på det medium, sätt och sammanhang i vilket Du Delar Bearbetningen.</li>
              <li id="s3b3" class="padding-left-normal padding-bottom-small">Du får inte erbjuda eller införa några ytterligare eller andra villkor eller tillämpa någon Teknisk skyddsåtgärd för Bearbetningar som begränsar nyttjandet av de rättigheter som ges enligt den Bearbetningslicens som Du tillämpar.</li>
            </ol>
          </li>
        
      </ol>
    </div>

    <!-- Section 4. Sui Generis Database Rights. -->
    <div class="padding-bottom-larger">
      <p id="s4" class="body-bigger padding-bottom-normal"><strong>Avsnitt 4 – Sui Generis-rättigheter för Databaser.</strong></p>
      <p class="body-big padding-bottom-normal">När Licensrättigheterna inkluderar Sui Generis-rättigheter för Databaser gäller följande för din användning av Licensmaterialet:</p>
      <ol type="a" class="body-big padding-left-normal">
          <li id="s4a" class="padding-left-normal padding-bottom-normal">
          
            för undvikande av missförstånd: avsnitt <a href="#s2a1">2(a)(1)</a> ger Dig rätt att extrahera, återanvända, mångfaldiga och Dela hela eller en väsentlig del av innehållet i databasen;
            
          </li>
          <li id="s4b" class="padding-left-normal padding-bottom-normal">
            
              om Du inkluderar hela eller en väsentlig del av databasinnehållet i en databas där Du har egna Sui generis-rättigheter för databasen, då är den databas som Du har Sui generis-rättigheter till (men inte dess innehåll) att betrakta som en Bearbetning, även vid tillämpning av avsnitt <a href="#s3b">3(b)</a>; och
            
          </li>
          <li id="s4c" class="padding-left-normal padding-bottom-small">Du måste uppfylla villkoren i avsnitt <a href="#s3a">3(a)</a> om Du Delar hela eller en väsentlig del av innehållet i databasen.</li>
      </ol>

      <span class="body-big">För undvikande av missförstånd: detta avsnitt <a href="#s4">4</a> kompletterar och ersätter inte Dina skyldigheter enligt denna Publika Licens när Licensrättigheterna inkluderar annan Upphovsrätt eller Liknande rättigheter.</span>
    </div>

    <!-- Section 5. Disclaimer -->
    <div class="padding-bottom-larger">
      <p id="s5" class="body-bigger padding-bottom-normal"><strong>Avsnitt 5 - Friskrivning från utfästelser och begränsning av ansvar.</strong></p>
      <ol style="font-weight: bold;" type="a" class="body-big padding-left-normal">
        <li id="s5a" class="padding-left-normal padding-bottom-normal"><strong>Om inte Licensgivaren har åtagit sig något annat och i den mån det är möjligt, erbjuder Licenstagaren Licenslicensmaterialet som det är och i den form det har gjorts tillgängligt, och gör inga utfästelser eller garantier av något slag rörande Licensmaterialet, vare sig uttryckliga, underförstådda, lagstadgade eller andra. Detta inkluderar, utan begränsning, garantier för titel, försäljningsbarhet, lämplighet för ett visst ändamål, icke-intrångsgörande, frånvaro av latenta eller andra defekter, korrekthet, eller närvaron eller frånvaron av fel, oavsett dessa är kända eller möjliga att upptäcka.Vid tillfällen där totala friskrivningar av utfästelser eller delar av dem inte är tillåtna är det möjligt att denna friskrivning inte gäller Dig.</strong></li>
        <li id="s5b" class="padding-left-normal padding-bottom-small"><strong>Licensgivaren kommer i möjligaste mån under inga omständigheter att ha något ansvar mot Dig på grund av någon rättsteori (inklusive, men utan begränsning, försumlighet) eller på annat sätt för några direkta, speciella, indirekta, tillfälliga, följdriktiga, straffrättsliga, exemplifierade eller andra förluster, kostnader , utgifter eller skador som följer av denna Publika Licens eller användning av Licensmaterialet, även om Licensgivaren har blivit upplyst om risken för sådana förluster, kostnader, utgifter eller skador. Vid tillfällen där en total ansvarsbegränsning eller en del av den inte är tillåten är det möjligt att denna begränsning inte gäller Dig.</strong></li>
      </ol>
      <ol start="3" type="a" class="body-big padding-left-normal">
        <li id="s5c" class="padding-left-normal padding-bottom-small">Den friskrivning från utfästelser och ansvarsbegränsning som anges ovan ska tolkas på ett sätt som, i den mån det är möjligt, mest liknar en absolut friskrivning och avstående från allt ansvar.</li>
      </ol>
    </div>

    <!-- Section 6. Term and Termination -->
    <div class="padding-bottom-larger">
      <p id="s6" class="body-bigger padding-bottom-normal"><strong>Avsnitt 6 – Giltighetstid och uppsägning.</strong></p>
      <ol type="a" class="body-big padding-left-normal">
        <li id="s6a" class="padding-left-normal padding-bottom-normal">Denna Publika Licens gäller under skyddstiden för den Upphovsrätt och/eller Liknande rättigheter som licensieras här. I den händelse Du underlåter att följa denna Publika Licens upphör dock automatiskt dina rättigheter enligt denna Publika Licens.</li>
        <li id="s6b" class="padding-left-normal padding-bottom-normal">
          <p class="body-big padding-bottom-normal">Om Din rätt att använda Licensmaterialet har upphört enligt 6(a), återinförs den:</p>
          <ol class="body-big padding-left-normal">
            <li id="s6b1" class="padding-left-normal padding-bottom-normal">automatiskt från den dag kränkningen upphörde, förutsatt att den upphörde inom 30 dagar från det att Du upptäckte kränkningen; eller</li>
            <li id="s6b2" class="padding-left-normal padding-bottom-small">vid uttryckligt återinförande av Licensgivaren.</li>
          </ol>
          För undvikande av missförstånd: detta avsnitt <a href="#s6b">6(b)</a> påverkar inte den rätt Licensgivaren kan ha att beivra Din kränkning av denna Publika Licens.
        </li>
        <li id="s6c" class="padding-left-normal padding-bottom-normal">För undvikande av missförstånd: Licensgivaren kan också erbjuda Licensmaterialet enligt separata villkor eller sluta distribuera Licensmaterialet när som helst; men att göra så innebär inte att denna Publika Licens upphör att gälla.</li>
        <li id="s6d" class="padding-left-normal padding-bottom-small">Avsnitten <a href="#s1">1</a>, <a href="#s5">5</a>, <a href="#s6">6</a>, <a href="#s7">7</a>, och <a href="#s8">8</a> gäller fortsatt även efter upphörandet av denna Publika Licens.</li>
      </ol>
    </div>

    <!-- Section 7. Other terms and conditions -->
    <div class="padding-bottom-larger">
      <p id="s7" class="body-bigger padding-bottom-normal"><strong>Avsnitt 7 – Övriga villkor.</strong></p>
      <ol type="a" class="body-big padding-left-normal">
        <li id="s7a" class="padding-left-normal padding-bottom-normal">Licensgivaren skall inte vara bunden av några ytterligare eller andra villkor som meddelats av Dig, om det inte uttryckligen överenskommits.</li>
        <li id="s7b" class="padding-left-normal padding-bottom-small">Alla överenskommelser, uppgörelser eller avtal om Licensmaterialet som inte anges här är skilda från och oberoende av villkoren i denna Publika Licens.</li>
      </ol>
    </div>

    <!-- Section 8. Interpretation -->
    <div class="padding-bottom-normal">
      <p id="s8" class="body-bigger padding-bottom-normal"><strong>Avsnitt 8 – Tolkning.</strong></p>
      <ol type="a" class="body-big padding-left-normal">
        <li id="s8a" class="padding-left-normal padding-bottom-normal">För undvikande av missförstånd: denna Publika Licens förminskar, avgränsar eller begränsar inte, och uppställer heller inte villkor för, någon användning av Licensmaterialet som lagligen kan företas utan tillstånd enligt denna Publika Licens, och ska heller inte tolkas så.</li>
        <li id="s8b" class="padding-left-normal padding-bottom-normal">Om någon bestämmelse i denna Publika Licens bedöms vara omöjlig att verkställa ska den i möjligaste mån automatiskt omvandlas i så liten utrsträckning som möjligt för att göra den verkställbar. Om bestämmelsen inte kan omvandlas ska den avskiljas från denna Publika Licens utan att påverka verkställigheten av de återstående villkoren.</li>
        <li id="s8c" class="padding-left-normal padding-bottom-normal">Inget villkor i denna Publika Licens ska avstås ifrån och ingen underlåtenhet att följa villkoren godkänns om inte Licensgivaren uttryckligen samtycker till det.</li>
        <li id="s8d" class="padding-left-normal">Ingenting i denna Publika Licens utgör eller får tolkas som en begränsning av eller avstående från några privilegier eller någon immunitet som Licensgivaren eller Du innehar, inklusive de som följer av rättspraxis hos någon domstol eller myndighet.</li>
      </ol>
    </div>
  </div>
</div>

<style>
  #legal-code-body {
    background-color: rgb(255, 255, 255);
    border: 5px solid rgb(176, 176, 176);
  }
</style>
  
      

<div id="legal-code-plain-text" style="font-weight: bold;" class="padding-vertical-normal" >
  <p class="body-big"><a href="#" class="link">View Legal Code as plain text</a></p>
</div>

      





<div id="about-cc-and-license" class="padding-bigger has-background-info-light" >
  <h4 class="padding-bottom-normal is-vcentered b-header"><i class="info icon padding-right-normal"></i>About Creative Commons</h4>
  <p class="has-text-black padding-left-big">
    Creative Commons is not a party to its public licenses. Notwithstanding, Creative Commons may elect to apply one of its public licenses to material it publishes and in those instances will be considered the "Licensor." The text of the Creative Commons public licenses is dedicated to the public domain under the <a href="#">CC0 Public Domain Dedication</a>. Except for the limited purpose of indicating that material is shared under a Creative Commons public license or as otherwise permitted by the Creative Commons policies published at <a href="creativecommons.org/policies">creativecommons.org/policies</a>, Creative Commons without its prior written consent including, without limitation, in connection with any unauthorized modifications to any of its public licenses or any other arrangements, understandings, or agreements concerning use of licensed material. For the avoidance of doubt, this paragraph does not form part of the public licenses.
  </p>
  <p class="has-text-black padding-left-big padding-top-normal">
    Creative Commons may be contacted at <a href="creativecommons.org">creativecommons.org</a>.
  </p>
</div>

      

<div
  class="menu padding-vertical-normal column is-half padding-right-large"
>
  <ul class="menu-list" >
    <li>
      
      
      
      
      <ul>
        
          <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="https://creativecommons.org/about/" class="is-inline body-big" style="font-weight: bold;">Learn more about our work</a></li>
        
        <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="https://creativecommons.org/about/cclicenses/" class="is-inline body-big" style="font-weight: bold;">Learn more about CC Licensing</a></li>
        <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="https://creativecommons.org/donate/" class="is-inline body-big" style="font-weight: bold;">Support our work</a></li>
        
          <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="https://chooser-beta.creativecommons.org/" class="is-inline body-big" style="font-weight: bold;">Use the license for your own material.<i class="icon external-link padding-bottom-small caption"></i></a></li>
        
      </ul>
    </li>
  </ul>
</div>

    </div>
  </div>

    </section>
  </main>
  
<footer class="main-footer margin-top-bigger">
  <div class="container">
    <div class="columns">
      <div class="column is-one-quarter">
        <a id="cc-footer-logo" href="https://creativecommons.org" class="main-logo margin-bottom-bigger has-text-white">
          <svg
  xmlns="http://www.w3.org/2000/svg"
  preserveAspectRatio="xMidYMid meet"
  viewBox="0 0 304 73">
  <use href="#logomark"></use>
  </svg></span>
        </a>
        <div>
          <address class="margin-bottom-normal">Creative Commons<br/>PO Box 1866, Mountain View CA 94042</address>
          <a href="mailto:info@creativecommons.org" class="mail">info@creativecommons.org</a><br/>
          <a href="tel://+1-415-429-6753" class="phone">+1-415-429-6753</a>
        </div>
        <div class="margin-vertical-large">
          <a href="https://www.instagram.com/creativecommons" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">instagram</i>
          </a>
          <a href="https://www.twitter.com/creativecommons" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">twitter</i>
          </a>
          <a href="https://www.facebook.com/creativecommons" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">facebook</i>
          </a>
          <a href="https://www.linkedin.com/company/creative-commons/" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">linkedin</i>
          </a>
        </div>
      </div>
      <div class="column is-three-quarters">
        <div class="columns">
          <div class="column is-full">
            <nav class="footer-navigation">
              <ul class="menu">
                <li><a href="#" class="menu-item">Who We Are</a></li>
                <li><a href="#" class="menu-item">What We Do</a></li>
                <li><a href="#" class="menu-item">Our Impact<i class="icon external-link"></i></a></li>
                <li><a href="#" class="menu-item">News</a></li>
              </ul>
            </nav>
          </div>
        </div>
        <div class="columns">
          <div class="column is-two-thirds">
            <div class="subscription">
              <h5 class="b-header">Subscribe to our newsletter</h5>
              <form class="newsletter">
                <input type="text" class="input" placeholder="Your email">
                <input type="submit" value="subscribe" class="button small">
              </form>
            </div>
            <div class="attribution margin-top-bigger">
              <p class="caption">
                Except where otherwise <a href="https://creativecommons.org/policies#license" target="_blank" rel="noopener">noted</a>, content on this site is licensed under a <a href="https://creativecommons.org/licenses/by/4.0/" target="_blank" rel="noopener">Creative Commons Attribution 4.0 International license</a>. <a href="https://creativecommons.org/website-icons" target="_blank" rel="noopener">Icons</a> by <a href="https://fontawesome.com/" target="_blank" rel="noopener">Font Awesome</a>.
              </p>
              <div class="margin-top-smaller">
                <i class="icon margin-right-small is-size-4">cclogo</i>
                <i class="icon margin-right-small is-size-4">ccby</i>
              </div>
            </div>
          </div>
          <div class="column is-one-third">
            <aside class="donate-section">
              <h5>Our work relies on you!</h5>
              <p>Help us keep the internet free and open.</p>
              <a class="button small donate" href="http://creativecommons.org/donate">
                <i class="icon cc-letterheart margin-right-small is-size-5 padding-top-smaller"></i>
                Donate now
              </a>
            </aside>
          </div>
        </div>
      </div>
    </div>
  </div>
  </footer>


  <script src="https://cdn.jsdelivr.net/npm/@creativecommons/vocabulary/js/vocabulary.js"></script>

  <script>
      /**
      * Get the fully-qualified URL of a Vocabulary asset.
      *
      * @param {string} version - the Vocabulary version in which to locate the asset
      * @param {string} path - the path of the asset being patched
      * @return {string} the fully qualified URL of the asset
      */
      const getFullyQualifiedUrl = (version, path) => {
      //   let baseUrl = 'https://unpkg.com/@creativecommons/vocabulary'
        // If you prefer jsDelivr instead, use
        let baseUrl = 'https://cdn.jsdelivr.net/npm/@creativecommons/vocabulary'
        return `${baseUrl}@${version}/${path}`
      }

      /**
      * Create an invisible container and place the asset into the DOM.
      *
      * This function is intended to be used to patch SVG assets that are later
      * referenced inside `<use>` tags in `<svg>` tags. It can also be used to force
      * an image to be downloaded to speed up its loading when referenced again.
      *
      * @param {string} path - the path of the asset being patched
      * @param {string} version - the Vocabulary version in which to locate the asset
      */
      const patchAssetIntoDom = (path, version = 'latest') => {
        fetch(getFullyQualifiedUrl(version, path)).then(response => {
          return response.text()
        }).then(data => {
          // Render SVG in the page
          const logo = document.querySelector('#cc-logo')
          const footerLogo = document.querySelector('#cc-footer-logo')
          logo.innerHTML = data;
          footerLogo.innerHTML = data;
        })
      }

      patchAssetIntoDom('assets/logos/cc/logomark.svg');

      /** Next Button On Click Event Listener **/
      document.getElementById("next-btn").addEventListener("click", function (e) {
        /**
        * On click redirect the user to page they are trying to visit
        * which is stored in the data-href.
        **/
        return window.location.href = this.dataset.href
      })
    </script>
    
  <script>
    /*
      Show/Hide Functionality for expand/collapse sections in use_of_licenses.html
    */
    let arrowArray = Array.from(document.getElementsByClassName("angle-down"))
    arrowArray.forEach(function(arrow) {
      arrow.addEventListener("click", handleArrowClicked);
    });

    function handleArrowClicked() {
      // Toggle consideration section's screen reader announcement text (inside of icon)
      if (this.dataset.consideration === "1" && this.dataset.direction === "down") {
        this.firstChild.innerHTML = "Hide Considerations for Licensors"
      } else if (this.dataset.consideration !== "1" && this.dataset.direction === "down") {
        this.firstChild.innerHTML = "Hide Considerations for the Public"
      } else if (this.dataset.consideration === "1" && this.dataset.direction === "up") {
        this.firstChild.innerHTML = "Show Considerations for Licensors"
      } else {
        this.firstChild.innerHTML = "Show Considerations for the Public"
      }
      // Toggle icon between up and down
      if (this.dataset.direction === "down") {
        // toggle icon to up arrow icon
        this.classList.remove("angle-down")
        this.classList.add("angle-up")
        this.dataset.direction = "up"
        // show <p> tag
        this.parentNode.parentNode.nextSibling.nextSibling.classList.remove("is-hidden");
      } else {
        // toggle icon to up arrow icon
        this.classList.add("angle-down")
        this.classList.remove("angle-up")
        this.dataset.direction = "down"
        // hide <p> tag
        this.parentNode.parentNode.nextSibling.nextSibling.classList.add("is-hidden");
      }
    };

  </script>

  </body>
</html>

<style>
body {
  background-color: rgb(245, 245, 245);
}

html[dir="rtl"] nav.breadcrumb>ul li+li:before {
  transform: scaleX(-1);
}

html[dir="rtl"] .breadcrumb li:first-child a {
    padding-right: 0;
    padding-left: .5rem;
}
</style>

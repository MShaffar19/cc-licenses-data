

<!DOCTYPE html>


<html lang="sv" class="no-js" dir="ltr">
<head about="http://creativecommons.org/licenses/by/4.0/">
    <meta charset="utf-8">
    <title>Creative Commons &mdash;  </title>
    <meta name="viewport" content="width=device-width, initial-scale=1.0">
    <meta name="description" content="">
    <meta name="author" content="">
    <meta http-equiv="Content-Type" content="application/xhtml+xml; charset=utf-8" />
    <meta name="keywords" content="">
    <link rel="stylesheet" href="https://cdn.jsdelivr.net/npm/bulma@0.9.0/css/bulma.min.css">
    <link rel="stylesheet" href="https://cdn.jsdelivr.net/npm/@creativecommons/vocabulary/css/vocabulary.css">
</head>
<body typeoff="cc:License">
  <style>svg { height: 73px; }</style>

<header>
  <nav class="navbar">
    <div class="navbar-brand">
      <a id="cc-logo" class="has-text-black" href="https://creativecommons.org" rel="home">
        <svg
          xmlns="http://www.w3.org/2000/svg"
          preserveAspectRatio="xMidYMid meet"
          viewBox="0 0 304 73">
        <!-- Automatically finds ID amongst all assets loaded using `patchAssetIntoDom()` -->
          <use href="#logomark"></use>
        </svg>
      </a>
      <a role="button" class="navbar-burger is-active" aria-label="menu" aria-expanded="false">
        <span aria-hidden="true"></span>
        <span aria-hidden="true"></span>
        <span aria-hidden="true"></span>
      </a>
    </div>
    <div class="navbar-menu is-active">
      <div class="navbar-end">
        <div class="navbar-item has-dropdown is-hoverable">
          <a class="navbar-link is-arrowless">Who We Are<i class="icon caret-down"></i></a>
          <div class="navbar-dropdown">
            <a class="navbar-item">Item 1</a>
            <a class="navbar-item">Item 2</a>
            <a class="navbar-item">Item 3</a>
          </div>
        </div>
        <div class="navbar-item has-dropdown is-hoverable">
          <a class="navbar-link is-arrowless">What We Do<i class="icon caret-down"></i></a>
          <div class="navbar-dropdown">
            <a class="navbar-item">Item 1</a>
            <a class="navbar-item">Item 2</a>
            <a class="navbar-item">Item 3</a>
          </div>
        </div>
        <a class="navbar-item">
          Our Impact<i class="icon external-link"></i>
        </a>
        <a class="navbar-item">
          News
        </a>
      </div>
    </div>
  </nav>
</header>

<style>
  html[dir="rtl"] .has-dropdown .navbar-link {
      flex-direction: row-reverse;
  }

  html[dir="rtl"] .navbar-end {
      margin-right: auto;
      margin-left: 0;
      justify-content: flex-start;
  }
</style>

  <main>
    <div class="level padding-left-big padding-right-large padding-vertical-normal">
          


<a class="skip-link" href="#content" >Hoppa över till innehåll</a>

<style>
  a.skip-link {
    left:-999px;
    position:absolute;
    top:auto;
    width:1px;
    height:1px;
    overflow:hidden;
    z-index:-999;
}
a.skip-link:focus, a.skip-link:active {
    color: black;
    font-weight: bolder;
    left: auto;
    top: auto;
    width: 30%;
    height: auto;
    overflow:auto;
    margin: 10px 35%;
    padding:5px;
    background-color: rgb(255, 255, 255);
    border-top: 10px solid rgb(60, 92, 153);
    border-bottom: 5px solid rgb(176, 176, 176);
    border-left: 5px solid rgb(176, 176, 176);
    border-right: 5px solid rgb(176, 176, 176);
    text-align:center;
    font-size:1.2em;
    z-index:999;
}
</style>

          <nav class="breadcrumb level-left caption bold" aria-label="breadcrumbs">
            <ul>
                <li><a href="#">Hem</a></li>
                <li><a href="#">License</a></li>
                <li class="is-active"><a href="#" aria-current="page displayed">
  License Deed for 


Erkännande 4.0 Internationell


</a></li>
            </ul>
          </nav>
          
            


<div class="locale level-right level-item has-text-black" >
  Languages available
  <div class="control margin-left-small">
    <div class="select">
      <select id="languages-dropdown">
        
        <option disabled>Select</option>

        
          <option
            id="option-id"
            
            value="id"
            data-link="/licenses/by/4.0/deed.id"
          >
            Bahasa Indonesia
          </option>
        
          <option
            id="option-eu"
            
            value="eu"
            data-link="/licenses/by/4.0/deed.eu"
          >
            Basque
          </option>
        
          <option
            id="option-de"
            
            value="de"
            data-link="/licenses/by/4.0/deed.de"
          >
            Deutsch
          </option>
        
          <option
            id="option-en"
            
            value="en"
            data-link="/licenses/by/4.0/"
          >
            English
          </option>
        
          <option
            id="option-es"
            
            value="es"
            data-link="/licenses/by/4.0/deed.es"
          >
            español
          </option>
        
          <option
            id="option-fr"
            
            value="fr"
            data-link="/licenses/by/4.0/deed.fr"
          >
            français
          </option>
        
          <option
            id="option-hr"
            
            value="hr"
            data-link="/licenses/by/4.0/deed.hr"
          >
            Hrvatski
          </option>
        
          <option
            id="option-it"
            
            value="it"
            data-link="/licenses/by/4.0/deed.it"
          >
            italiano
          </option>
        
          <option
            id="option-lv"
            
            value="lv"
            data-link="/licenses/by/4.0/deed.lv"
          >
            latviešu
          </option>
        
          <option
            id="option-lt"
            
            value="lt"
            data-link="/licenses/by/4.0/deed.lt"
          >
            Lietuviškai
          </option>
        
          <option
            id="option-mi"
            
            value="mi"
            data-link="/licenses/by/4.0/deed.mi"
          >
            Māori
          </option>
        
          <option
            id="option-nl"
            
            value="nl"
            data-link="/licenses/by/4.0/deed.nl"
          >
            Nederlands
          </option>
        
          <option
            id="option-no"
            
            value="no"
            data-link="/licenses/by/4.0/deed.no"
          >
            norsk
          </option>
        
          <option
            id="option-pl"
            
            value="pl"
            data-link="/licenses/by/4.0/deed.pl"
          >
            polski
          </option>
        
          <option
            id="option-pt"
            
            value="pt"
            data-link="/licenses/by/4.0/deed.pt"
          >
            Português
          </option>
        
          <option
            id="option-ro"
            
            value="ro"
            data-link="/licenses/by/4.0/deed.ro"
          >
            Română
          </option>
        
          <option
            id="option-sl"
            
            value="sl"
            data-link="/licenses/by/4.0/deed.sl"
          >
            Slovenščina
          </option>
        
          <option
            id="option-fi"
            
            value="fi"
            data-link="/licenses/by/4.0/deed.fi"
          >
            suomi
          </option>
        
          <option
            id="option-sv"
            selected
            value="sv"
            data-link="/licenses/by/4.0/deed.sv"
          >
            svenska
          </option>
        
          <option
            id="option-tr"
            
            value="tr"
            data-link="/licenses/by/4.0/deed.tr"
          >
            Türkçe
          </option>
        
          <option
            id="option-cs"
            
            value="cs"
            data-link="/licenses/by/4.0/deed.cs"
          >
            česky
          </option>
        
          <option
            id="option-el"
            
            value="el"
            data-link="/licenses/by/4.0/deed.el"
          >
            Ελληνικά
          </option>
        
          <option
            id="option-ru"
            
            value="ru"
            data-link="/licenses/by/4.0/deed.ru"
          >
            Русский
          </option>
        
          <option
            id="option-uk"
            
            value="uk"
            data-link="/licenses/by/4.0/deed.uk"
          >
            Українська
          </option>
        
          <option
            id="option-ar"
            
            value="ar"
            data-link="/licenses/by/4.0/deed.ar"
          >
            العربيّة
          </option>
        
          <option
            id="option-ja"
            
            value="ja"
            data-link="/licenses/by/4.0/deed.ja"
          >
            日本語
          </option>
        
          <option
            id="option-zh-Hans"
            
            value="zh-Hans"
            data-link="/licenses/by/4.0/deed.zh-Hans"
          >
            简体中文
          </option>
        
          <option
            id="option-zh-Hant"
            
            value="zh-Hant"
            data-link="/licenses/by/4.0/deed.zh-Hant"
          >
            繁體中文
          </option>
        
          <option
            id="option-ko"
            
            value="ko"
            data-link="/licenses/by/4.0/deed.ko"
          >
            한국어
          </option>
        

        
      </select>
    </div>
    <div class="icon is-small is-left">
      <!-- TODO Add icons here -->
    </div>
  </div>
</div>

<script>
  const select = document.getElementById("languages-dropdown")

  select.addEventListener("input", function () {
    const language_code = select.value
    const option = document.getElementById("option-" + language_code)
    window.location.href = option.dataset.link
  })
</script>

          
    </div>
    <section id="content" class="padding-horizontal-larger">
      
<div class="level container">
  <div class="level-item level-right">
    <button id="next-btn" class="button tiny is-pulled-right" data-href="/licenses/by/4.0/legalcode.sv">See the legal code</button>
  </div>
</div>

      
  <div class="container">
    
<div id="deed-body" class="margin-vertical-bigger padding-xxl" >
  

<h3 class="is-vcentered is-hidden-touch">
  
    <span class="padding-right-bigger">
    
      





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


    </span>
  CC BY 4.0
</h3>
<h3 class="is-vcentered is-hidden-desktop is-hidden-mobile has-text-centered">
  
    <span class="padding-right-big">
    
      





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


      





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small"
></i>


    </span>
    CC BY 4.0
</h3>
<h3 class="is-hidden-tablet has-text-centered">
  
    <span>
    
      





<i
  class="cc-logo icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-logo icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


      





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


      





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


      





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch margin-normal padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop margin-small padding-bottom-small margin-horizontal-smaller margin-vertical-small"
></i>


    </span>
</h3>
<h4 class="has-text-centered is-hidden-tablet padding-left-normal">CC BY 4.0</h4>
<h2 class="margin-bottom-larger b-header is-hidden-touch">


Erkännande 4.0 Internationell

</h2>
<h3 class="margin-bottom-larger b-header is-hidden-desktop has-text-centered">


Erkännande 4.0 Internationell

</h3>

  
  
  <h3 class="b-header has-text-black padding-bottom-big padding-top-normal" style="font-weight: bold;">Du har tillstånd att:</h3>
  <p class="has-text-black body-big padding-bottom-normal"><strong>Dela</strong> &mdash; kopiera och vidaredistribuera materialet oavsett medium eller format
  </p>
  <p class="has-text-black body-big padding-bottom-small"><strong>Bearbeta</strong> &mdash; remixa, transformera, och bygg vidare på materialet
  </p>
  <p class="has-text-black body-big padding-bottom-small">
    Licensgivaren kan inte återkalla dessa friheter så länge du följer licensvillkoren.
  </p>
  <h3 class="b-header has-text-black padding-bottom-big padding-top-normal" style="font-weight: bold;">
    På följande villkor:
  </h3>
  <div class="columns is-multiline">
    
    <div class="column is-1">
      





<i
  class="cc-by icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch "
></i>
<i
  class="cc-by icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop "
></i>


    </div>
    <div class="column is-11">
      <p class="has-text-black body-big padding-bottom-normal">
        <span style="font-weight: bold;">Erkännande</span> -

        Du måste ge <a href="#" id="appropriate_credit_popup" class="helpLink">ett korrekt erkännande</a></span>, ange en hyperlänk till licensen, och <span rel="cc:requires" resource="http://creativecommons.org/ns#Notice"><a href="#" id="indicate_changes_popup" class="helpLink">ange om bearbetningar är gjorda </a></span>.  Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att licensgivaren stödjer dig eller ditt användande.
      </p>
    </div>
    
    <div class="column is-1">
      





<i
  class="cc-nc icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch "
></i>
<i
  class="cc-nc icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop "
></i>


    </div>
    <div class="column is-11">
      <p class="has-text-black body-big padding-bottom-normal">
        <span style="font-weight: bold;">IckeKommersiell</span> -

        Du får inte använda materialet för <a href="#" id="commercial_purposes_popup" class="helpLink">kommersiella ändamål</a>.
      </p>
    </div>
    <div class="column is-1">
      





<i
  class="cc-sa icon has-text-black has-background-white is-size-1 padding-left-big is-hidden-touch "
></i>
<i
  class="cc-sa icon has-text-black has-background-white is-size-2 padding-left-normal is-hidden-desktop "
></i>


    </div>
    <div class="column is-11">
      <p class="has-text-black body-big padding-bottom-normal">
        <span style="font-weight: bold;">DelaLika</span> - Om du remixar, transformerar eller bygger vidare på materialet måste du distribuera dina bidrag under <a href="#" id="same_license_popup" class="helpLink">samma licens</a> som originalet.
      </p>
    </div>
    <div class="column is-1">
    </div>
    <div class="column is-11">
      <p class="has-text-black body-big padding-bottom-normal">
        <span style="font-weight: bold;">Inga ytterligare begränsningar</span> - Du får inte tillämpa lagliga begränsningar eller <a href="#" id="technological_measures_popup" class="helpLink">teknologiska metoder</a> som juridiskt begränsar andra från att gör något som licensen tillåter. 
      </p>
    </div>
  </div>
  <h3 class="b-header has-text-black padding-bottom-big padding-top-normal" style="font-weight: bold;">Anmärkningar:</h3>
  <p class="has-text-black body-big padding-bottom-normal">
    Du behöver inte följa licensvillkoren för de delar av materialet som finns i public domain eller där ditt användande är tillåtet av en tillämplig <a href="#" id="exception_or_limitation_popup" class="helpLink">undantag eller begränsning</a>.
  </p>
  <p class="has-text-black body-big padding-bottom-normal">
    Inga garantier ges. Licensen ger eller ger dig inte alla de nödvändiga villkoren för ditt tänkta användande av verket. Till exempel, andra rättigheter som <a href="#" id="publicity_privacy_or_moral_rights_popup" class="helpLink">publicitet, integritetslagstiftning, eller ideella rättigheter </a> kan begränsa hur du kan använda verket. 
  </p>
</div>

<style>
  #deed-body {
    background-color: rgb(255, 255, 255);
    border-top: 10px solid rgb(60, 92, 153);
    border-bottom: 5px solid rgb(176, 176, 176);
    border-left: 5px solid rgb(176, 176, 176);
    border-right: 5px solid rgb(176, 176, 176);
  }
</style>

    






<div id="disclaimer-info-section" class="padding-bigger has-background-info-light" >
  <h4 class="padding-bottom-normal is-vcentered b-header"><i class="info icon padding-right-normal"></i>Friskrivning</h4>
  <p class="has-text-black padding-left-big">
    Denna sammanfattning uppmärksammar enbart vissa av de viktigaste inslagen och villkoren från den faktiska licensen. Den är inte en licens och har inget juridiskt värde. Du bör noggrant gå igenom alla villkor i den faktiska licensen innan du använder det licensierade materialet.
  </p>
  <p class="has-text-black padding-left-big padding-top-normal">
    Creative Commons är ingen advokatbyrå och tillhandahåller inga juridiska tjänster eller juridisk rådgivning. Distribution eller visning av, samt länkning till denna handling eller licensen som sammanfattas skapar ingen advokat-klient- eller annat förhållande.
  </p>
</div>

    <div class="columns margin-top-normal is-vcentered" >
      

<div
  class="menu padding-vertical-normal column is-half padding-right-large"
>
  <ul class="menu-list" >
    <li>
      
      
      
        <p class="body-big has-text-black">
          Creative Commons is the nonprofit behind the open licenses that allow creators to share their work. Our licenses and legal tools are free to use.
        </p>
      
      
      <ul>
        
          <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="#" class="is-inline body-big" style="font-weight: bold;">Learn more about our work</a></li>
        
        <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="#" class="is-inline body-big" style="font-weight: bold;">Learn more about CC Licensing</a></li>
        <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="#" class="is-inline body-big" style="font-weight: bold;">Support our work</a></li>
        
          <li><span class="body-bigger padding-right-normal padding-top-small">&#8226;</span><a href="#" class="is-inline body-big" style="font-weight: bold;">Use the license for your own material.<i class="icon external-link padding-bottom-small caption"></i></a></li>
        
      </ul>
    </li>
  </ul>
</div>

      

<div
  id="column is-full margin-top-bigger"
  style="width: 100%;"

>
  <div class="card entry-post">
    <div class="card-content">
      <h4>Get The Latest Updates</h4>
      <p class="body-big">Subscribe to our monthly newsletter.</p>
      <form class="margin-top-normal">
        <div class="field has-addons">
          <label for="email" class="is-sr-only">Email address</label>
          <input type="text" id="email" class="input is-medium" placeholder="Email Address">
          <button type="submit" class="button is-primary">Join</button>
        </div>
      </form>
    </div>
  </div>
</div>

    </div>
  </div>

    </section>
  </main>
  
<footer class="main-footer margin-top-bigger">
  <div class="container">
    <div class="columns">
      <div class="column is-one-quarter">
        <a id="cc-footer-logo" href="https://creativecommons.org" class="main-logo margin-bottom-bigger has-text-white">
          <svg
  xmlns="http://www.w3.org/2000/svg"
  preserveAspectRatio="xMidYMid meet"
  viewBox="0 0 304 73">
  <use href="#logomark"></use>
  </svg></span>
        </a>
        <div>
          <address class="margin-bottom-normal">Creative Commons<br/>PO Box 1866, Mountain View CA 94042</address>
          <a href="mailto:info@creativecommons.org" class="mail">info@creativecommons.org</a><br/>
          <a href="tel://+1-415-429-6753" class="phone">+1-415-429-6753</a>
        </div>
        <div class="margin-vertical-large">
          <a href="https://www.instagram.com/creativecommons" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">instagram</i>
          </a>
          <a href="https://www.twitter.com/creativecommons" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">twitter</i>
          </a>
          <a href="https://www.facebook.com/creativecommons" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">facebook</i>
          </a>
          <a href="https://www.linkedin.com/company/creative-commons/" class="social has-text-white" target="_blank" rel="noopener">
            <i class="icon margin-right-small is-size-4">linkedin</i>
          </a>
        </div>
      </div>
      <div class="column is-three-quarters">
        <div class="columns">
          <div class="column is-full">
            <nav class="footer-navigation">
              <ul class="menu">
                <li><a href="#" class="menu-item">Who We Are</a></li>
                <li><a href="#" class="menu-item">What We Do</a></li>
                <li><a href="#" class="menu-item">Our Impact<i class="icon external-link"></i></a></li>
                <li><a href="#" class="menu-item">News</a></li>
              </ul>
            </nav>
          </div>
        </div>
        <div class="columns">
          <div class="column is-two-thirds">
            <div class="subscription">
              <h5 class="b-header">Subscribe to our newsletter</h5>
              <form class="newsletter">
                <input type="text" class="input" placeholder="Your email">
                <input type="submit" value="subscribe" class="button small">
              </form>
            </div>
            <div class="attribution margin-top-bigger">
              <p class="caption">
                Except where otherwise <a href="https://creativecommons.org/policies#license" target="_blank" rel="noopener">noted</a>, content on this site is licensed under a <a href="https://creativecommons.org/licenses/by/4.0/" target="_blank" rel="noopener">Creative Commons Attribution 4.0 International license</a>. <a href="https://creativecommons.org/website-icons" target="_blank" rel="noopener">Icons</a> by <a href="https://fontawesome.com/" target="_blank" rel="noopener">Font Awesome</a>.
              </p>
              <div class="margin-top-smaller">
                <i class="icon margin-right-small is-size-4">cclogo</i>
                <i class="icon margin-right-small is-size-4">ccby</i>
              </div>
            </div>
          </div>
          <div class="column is-one-third">
            <aside class="donate-section">
              <h5>Our work relies on you!</h5>
              <p>Help us keep the internet free and open.</p>
              <a class="button small donate" href="http://creativecommons.org/donate">
                <i class="icon cc-letterheart margin-right-small is-size-5 padding-top-smaller"></i>
                Donate now
              </a>
            </aside>
          </div>
        </div>
      </div>
    </div>
  </div>
  </footer>


  <script src="https://cdn.jsdelivr.net/npm/@creativecommons/vocabulary/js/vocabulary.js"></script>

  <script>
      /**
      * Get the fully-qualified URL of a Vocabulary asset.
      *
      * @param {string} version - the Vocabulary version in which to locate the asset
      * @param {string} path - the path of the asset being patched
      * @return {string} the fully qualified URL of the asset
      */
      const getFullyQualifiedUrl = (version, path) => {
      //   let baseUrl = 'https://unpkg.com/@creativecommons/vocabulary'
        // If you prefer jsDelivr instead, use
        let baseUrl = 'https://cdn.jsdelivr.net/npm/@creativecommons/vocabulary'
        return `${baseUrl}@${version}/${path}`
      }

      /**
      * Create an invisible container and place the asset into the DOM.
      *
      * This function is intended to be used to patch SVG assets that are later
      * referenced inside `<use>` tags in `<svg>` tags. It can also be used to force
      * an image to be downloaded to speed up its loading when referenced again.
      *
      * @param {string} path - the path of the asset being patched
      * @param {string} version - the Vocabulary version in which to locate the asset
      */
      const patchAssetIntoDom = (path, version = 'latest') => {
        fetch(getFullyQualifiedUrl(version, path)).then(response => {
          return response.text()
        }).then(data => {
          // Render SVG in the page
          const logo = document.querySelector('#cc-logo')
          const footerLogo = document.querySelector('#cc-footer-logo')
          logo.innerHTML = data;
          footerLogo.innerHTML = data;
        })
      }

      patchAssetIntoDom('assets/logos/cc/logomark.svg');

      /** Next Button On Click Event Listener **/
      document.getElementById("next-btn").addEventListener("click", function (e) {
        /**
        * On click redirect the user to page they are trying to visit
        * which is stored in the data-href.
        **/
        return window.location.href = this.dataset.href
      })
    </script>
    
    
  </body>
</html>

<style>
body {
  background-color: rgb(245, 245, 245);
}

html[dir="rtl"] nav.breadcrumb>ul li+li:before {
  transform: scaleX(-1);
}

html[dir="rtl"] .breadcrumb li:first-child a {
    padding-right: 0;
    padding-left: .5rem;
}
</style>
